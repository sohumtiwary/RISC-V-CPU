module scoreboard;
  // For Milestone 0, we’ll just check final reg values in tb_top.
  // This file stays as a placeholder for later (ISA-model scoreboard).
endmodule
